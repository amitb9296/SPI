module tb_spi;
	reg 		 clk,    // Clock
	reg 		 rst,    // Asynchronous reset active high
	reg  [7:0]   din,dvsr,
	reg 		 wr,
	wire [7:0]   dout,
	wire         spi_clk,spi_mosi,
	reg          spi_miso,
	wire         spi_done, spi_idle



endmodule